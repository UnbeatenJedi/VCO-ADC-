//Verilog HDL for "vco_adc", "digi_inv" "functional"


module digi_inv (input x, output y );
assign y = !x;

endmodule

//Verilog HDL for "vco_adc", "inverter" "functional"


module inverter ( );

endmodule

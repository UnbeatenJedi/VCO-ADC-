//Verilog HDL for "vco_adc", "inverter23" "functional"


module inverter23 ( );

endmodule
